--------------------------------------------------------------------------------
-- File: basic_app_types_pkg.vhd
-- Author: Stub package for P2 FSM compilation test
-- Date: 2025-11-05
-- Version: 0.1 (STUB)
--
-- Description:
--   Minimal stub package for basic_app_types_pkg.
--   Provides type definitions for Basic Probe Driver application.
--
-- Status: STUB - Will be replaced by forge-codegen generated code
--
-- Note: This is a minimal stub to satisfy dependency checking during
--       initial FSM compilation. The real package will be generated from
--       basic_probe_driver.yaml using forge-codegen tools.
--------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package basic_app_types_pkg is

    ----------------------------------------------------------------------------
    -- Basic Data Types
    --
    -- TODO: Add application-specific types here when generated from YAML
    ----------------------------------------------------------------------------

    -- Placeholder: No types currently required by FSM
    -- The FSM uses standard IEEE types (std_logic, unsigned, signed)

end package basic_app_types_pkg;

package body basic_app_types_pkg is

    -- No functions or procedures yet

end package body basic_app_types_pkg;
