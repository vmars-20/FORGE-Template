--------------------------------------------------------------------------------
-- File: basic_app_voltage_pkg.vhd
-- Author: Stub package for P2 FSM compilation test
-- Date: 2025-11-05
-- Version: 0.1 (STUB)
--
-- Description:
--   Minimal stub package for basic_app_voltage_pkg.
--   Provides voltage conversion utilities for Basic Probe Driver.
--
-- Status: STUB - Will be replaced by forge-codegen generated code
--
-- Note: This is a minimal stub to satisfy dependency checking during
--       initial FSM compilation. The real package will be generated from
--       basic_probe_driver.yaml using forge-codegen tools.
--------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package basic_app_voltage_pkg is

    ----------------------------------------------------------------------------
    -- Voltage Conversion Functions
    --
    -- TODO: Add voltage conversion functions when generated from YAML:
    --   - mV_to_dac_code()
    --   - dac_code_to_mV()
    --   - voltage range constants
    ----------------------------------------------------------------------------

    -- Placeholder: No voltage functions currently called by FSM

end package basic_app_voltage_pkg;

package body basic_app_voltage_pkg is

    -- No functions or procedures yet

end package body basic_app_voltage_pkg;
